//----------------------------------------------------------------
// SoC Buttom interface behavioural
// Support: Debounce
// Last Modified Date: 2023/7/17
// Version: 1.0
// Author: Clark Pu
//----------------------------------------------------------------


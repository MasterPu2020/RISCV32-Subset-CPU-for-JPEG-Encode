//----------------------------------------------------------------
// Asynchronous single port read-only memory behavioural
// Support: 32-bit read, address add by 4
// Last Modified Date: 2023/7/17
// Version: 1.0
// Author: Clark Pu
//----------------------------------------------------------------

module rom #(parameter WIDTH = 32, DEPTH = 2048) (
  input wire [WIDTH-1:0] address,
  output wire [WIDTH-1:0] rdata
);

  wire [WIDTH-1:0] memory [DEPTH-1:0];
  assign rdata = memory[address[WIDTH-1:2]];

  // JPEG encode program
  assign memory[   0] = 32'h00005093;
  assign memory[   1] = 32'h0FA05113;
  assign memory[   2] = 32'h01005193;
  assign memory[   3] = 32'h00005213;
  assign memory[   4] = 32'h00B05293;
  assign memory[   5] = 32'h01005313;
  assign memory[   6] = 32'h04114463;
  assign memory[   7] = 32'h1000A9A3;
  assign memory[   8] = 32'h3200A0A3;
  assign memory[   9] = 32'h00105393;
  assign memory[  10] = 32'h0053DC63;
  assign memory[  11] = 32'h00138433;
  assign memory[  12] = 32'h103429A3;
  assign memory[  13] = 32'h323420A3;
  assign memory[  14] = 32'h0013D393;
  assign memory[  15] = 32'hFE0006E3;
  assign memory[  16] = 32'h0063DC63;
  assign memory[  17] = 32'h00138433;
  assign memory[  18] = 32'h100429A3;
  assign memory[  19] = 32'h320420A3;
  assign memory[  20] = 32'h0013D393;
  assign memory[  21] = 32'hFE0006E3;
  assign memory[  22] = 32'h0100D093;
  assign memory[  23] = 32'hFA000EE3;
  assign memory[  24] = 32'h41C05093;
  assign memory[  25] = 32'h49B05113;
  assign memory[  26] = 32'h02005F13;
  assign memory[  27] = 32'h00B05F93;
  assign memory[  28] = 32'h01FF1F33;
  assign memory[  29] = 32'h00005F93;
  assign memory[  30] = 32'h01FF61B3;
  assign memory[  31] = 32'h00114863;
  assign memory[  32] = 32'h0030A023;
  assign memory[  33] = 32'h0010D093;
  assign memory[  34] = 32'hFE000AE3;
  assign memory[  35] = 32'h01605F93;
  assign memory[  36] = 32'hF4305E93;
  assign memory[  37] = 32'h01FE9EB3;
  assign memory[  38] = 32'h00B05F93;
  assign memory[  39] = 32'h4AC05F13;
  assign memory[  40] = 32'h01FF1F33;
  assign memory[  41] = 32'h01DF6EB3;
  assign memory[  42] = 32'h04205F93;
  assign memory[  43] = 32'h01DFE0B3;
  assign memory[  44] = 32'h4A102F23;
  assign memory[  45] = 32'h01605F93;
  assign memory[  46] = 32'hF6B05E93;
  assign memory[  47] = 32'h01FE9EB3;
  assign memory[  48] = 32'h00B05F93;
  assign memory[  49] = 32'h01005F13;
  assign memory[  50] = 32'h01FF1F33;
  assign memory[  51] = 32'h01DF6EB3;
  assign memory[  52] = 32'h31305F93;
  assign memory[  53] = 32'h01DFE133;
  assign memory[  54] = 32'h4A202E23;
  assign memory[  55] = 32'h01605F93;
  assign memory[  56] = 32'hFB405E93;
  assign memory[  57] = 32'h01FE9EB3;
  assign memory[  58] = 32'h00B05F93;
  assign memory[  59] = 32'h1CA05F13;
  assign memory[  60] = 32'h01FF1F33;
  assign memory[  61] = 32'h01DF6EB3;
  assign memory[  62] = 32'h60505F93;
  assign memory[  63] = 32'h01DFE1B3;
  assign memory[  64] = 32'h4A302DA3;
  assign memory[  65] = 32'h01605F93;
  assign memory[  66] = 32'hFDB05E93;
  assign memory[  67] = 32'h01FE9EB3;
  assign memory[  68] = 32'h00B05F93;
  assign memory[  69] = 32'h52F05F13;
  assign memory[  70] = 32'h01FF1F33;
  assign memory[  71] = 32'h01DF6EB3;
  assign memory[  72] = 32'h0D505F93;
  assign memory[  73] = 32'h01DFE233;
  assign memory[  74] = 32'h4A402FA3;
  assign memory[  75] = 32'h00105293;
  assign memory[  76] = 32'h00502D23;
  assign memory[  77] = 32'h205027A3;
  assign memory[  78] = 32'h225023A3;
  assign memory[  79] = 32'h00205313;
  assign memory[  80] = 32'h006020A3;
  assign memory[  81] = 32'h00602623;
  assign memory[  82] = 32'h10602A23;
  assign memory[  83] = 32'h10602AA3;
  assign memory[  84] = 32'h20602823;
  assign memory[  85] = 32'h20602D23;
  assign memory[  86] = 32'h20602DA3;
  assign memory[  87] = 32'h20602E23;
  assign memory[  88] = 32'h326020A3;
  assign memory[  89] = 32'h32602123;
  assign memory[  90] = 32'h00305393;
  assign memory[  91] = 32'h00702123;
  assign memory[  92] = 32'h007026A3;
  assign memory[  93] = 32'h00702723;
  assign memory[  94] = 32'h007027A3;
  assign memory[  95] = 32'h00702823;
  assign memory[  96] = 32'h007028A3;
  assign memory[  97] = 32'h10702B23;
  assign memory[  98] = 32'h20702EA3;
  assign memory[  99] = 32'h327021A3;
  assign memory[ 100] = 32'h00405413;
  assign memory[ 101] = 32'h008021A3;
  assign memory[ 102] = 32'h00802923;
  assign memory[ 103] = 32'h00802DA3;
  assign memory[ 104] = 32'h108029A3;
  assign memory[ 105] = 32'h10802BA3;
  assign memory[ 106] = 32'h12802223;
  assign memory[ 107] = 32'h20802F23;
  assign memory[ 108] = 32'h22802423;
  assign memory[ 109] = 32'h32802223;
  assign memory[ 110] = 32'h32802923;
  assign memory[ 111] = 32'h00505493;
  assign memory[ 112] = 32'h00902223;
  assign memory[ 113] = 32'h009029A3;
  assign memory[ 114] = 32'h10902C23;
  assign memory[ 115] = 32'h129022A3;
  assign memory[ 116] = 32'h12902A23;
  assign memory[ 117] = 32'h20902FA3;
  assign memory[ 118] = 32'h329022A3;
  assign memory[ 119] = 32'h32902323;
  assign memory[ 120] = 32'h34902123;
  assign memory[ 121] = 32'h34902923;
  assign memory[ 122] = 32'h00605513;
  assign memory[ 123] = 32'h00A022A3;
  assign memory[ 124] = 32'h00A02A23;
  assign memory[ 125] = 32'h14A02223;
  assign memory[ 126] = 32'h14A02A23;
  assign memory[ 127] = 32'h20A028A3;
  assign memory[ 128] = 32'h22A02023;
  assign memory[ 129] = 32'h32A023A3;
  assign memory[ 130] = 32'h32A029A3;
  assign memory[ 131] = 32'h36A02123;
  assign memory[ 132] = 32'h36A02923;
  assign memory[ 133] = 32'h00705593;
  assign memory[ 134] = 32'h00B02AA3;
  assign memory[ 135] = 32'h10B02CA3;
  assign memory[ 136] = 32'h12B02323;
  assign memory[ 137] = 32'h16B02223;
  assign memory[ 138] = 32'h16B02A23;
  assign memory[ 139] = 32'h22B020A3;
  assign memory[ 140] = 32'h32B02423;
  assign memory[ 141] = 32'h38B02123;
  assign memory[ 142] = 32'h38B02923;
  assign memory[ 143] = 32'h00805613;
  assign memory[ 144] = 32'h00C02B23;
  assign memory[ 145] = 32'h10C02D23;
  assign memory[ 146] = 32'h12C02AA3;
  assign memory[ 147] = 32'h18C02223;
  assign memory[ 148] = 32'h22C02123;
  assign memory[ 149] = 32'h32C02A23;
  assign memory[ 150] = 32'h34C021A3;
  assign memory[ 151] = 32'h34C029A3;
  assign memory[ 152] = 32'h3AC02123;
  assign memory[ 153] = 32'h00905693;
  assign memory[ 154] = 32'h00D02BA3;
  assign memory[ 155] = 32'h12D023A3;
  assign memory[ 156] = 32'h14D022A3;
  assign memory[ 157] = 32'h18D02A23;
  assign memory[ 158] = 32'h1AD02223;
  assign memory[ 159] = 32'h1AD02A23;
  assign memory[ 160] = 32'h22D021A3;
  assign memory[ 161] = 32'h32D024A3;
  assign memory[ 162] = 32'h32D02AA3;
  assign memory[ 163] = 32'h36D021A3;
  assign memory[ 164] = 32'h3AD02923;
  assign memory[ 165] = 32'h3CD02123;
  assign memory[ 166] = 32'h3CD02923;
  assign memory[ 167] = 32'h3ED02123;
  assign memory[ 168] = 32'h00A05713;
  assign memory[ 169] = 32'h00E02C23;
  assign memory[ 170] = 32'h10E02DA3;
  assign memory[ 171] = 32'h12E02B23;
  assign memory[ 172] = 32'h14E02AA3;
  assign memory[ 173] = 32'h1CE02223;
  assign memory[ 174] = 32'h1CE02A23;
  assign memory[ 175] = 32'h22E02223;
  assign memory[ 176] = 32'h22E024A3;
  assign memory[ 177] = 32'h32E02523;
  assign memory[ 178] = 32'h34E02223;
  assign memory[ 179] = 32'h34E02A23;
  assign memory[ 180] = 32'h36E029A3;
  assign memory[ 181] = 32'h40E028A3;
  assign memory[ 182] = 32'h00B05793;
  assign memory[ 183] = 32'h00F02E23;
  assign memory[ 184] = 32'h12F02423;
  assign memory[ 185] = 32'h16F022A3;
  assign memory[ 186] = 32'h1EF02223;
  assign memory[ 187] = 32'h20F021A3;
  assign memory[ 188] = 32'h22F022A3;
  assign memory[ 189] = 32'h22F02BA3;
  assign memory[ 190] = 32'h32F02B23;
  assign memory[ 191] = 32'h38F021A3;
  assign memory[ 192] = 32'h38F029A3;
  assign memory[ 193] = 32'h3EF02923;
  assign memory[ 194] = 32'h00C05813;
  assign memory[ 195] = 32'h030024A3;
  assign memory[ 196] = 32'h13002BA3;
  assign memory[ 197] = 32'h15002323;
  assign memory[ 198] = 32'h17002AA3;
  assign memory[ 199] = 32'h190022A3;
  assign memory[ 200] = 32'h330025A3;
  assign memory[ 201] = 32'h33002BA3;
  assign memory[ 202] = 32'h350022A3;
  assign memory[ 203] = 32'h35002AA3;
  assign memory[ 204] = 32'h00E05893;
  assign memory[ 205] = 32'h01102323;
  assign memory[ 206] = 32'h21102923;
  assign memory[ 207] = 32'h41102123;
  assign memory[ 208] = 32'h00F05913;
  assign memory[ 209] = 32'h19202AA3;
  assign memory[ 210] = 32'h35202323;
  assign memory[ 211] = 32'h41202923;
  assign memory[ 212] = 32'h01805993;
  assign memory[ 213] = 32'h23302523;
  assign memory[ 214] = 32'h01905A13;
  assign memory[ 215] = 32'h234025A3;
  assign memory[ 216] = 32'h01A05A93;
  assign memory[ 217] = 32'h01502EA3;
  assign memory[ 218] = 32'h255023A3;
  assign memory[ 219] = 32'h01B05B13;
  assign memory[ 220] = 32'h03602523;
  assign memory[ 221] = 32'h25602BA3;
  assign memory[ 222] = 32'h01C05B93;
  assign memory[ 223] = 32'h03702CA3;
  assign memory[ 224] = 32'h01E05C13;
  assign memory[ 225] = 32'h018023A3;
  assign memory[ 226] = 32'h218029A3;
  assign memory[ 227] = 32'h03805C93;
  assign memory[ 228] = 32'h23902623;
  assign memory[ 229] = 32'h03905D13;
  assign memory[ 230] = 32'h23A02C23;
  assign memory[ 231] = 32'h03A05D93;
  assign memory[ 232] = 32'h05B024A3;
  assign memory[ 233] = 32'h27B023A3;
  assign memory[ 234] = 32'h03B05E13;
  assign memory[ 235] = 32'h05C02CA3;
  assign memory[ 236] = 32'h27C02BA3;
  assign memory[ 237] = 32'h03E05E93;
  assign memory[ 238] = 32'h01D02423;
  assign memory[ 239] = 32'h21D02A23;
  assign memory[ 240] = 32'h07805093;
  assign memory[ 241] = 32'h00102F23;
  assign memory[ 242] = 32'h221026A3;
  assign memory[ 243] = 32'h07905113;
  assign memory[ 244] = 32'h022025A3;
  assign memory[ 245] = 32'h282023A3;
  assign memory[ 246] = 32'h07A05193;
  assign memory[ 247] = 32'h063024A3;
  assign memory[ 248] = 32'h28302BA3;
  assign memory[ 249] = 32'h07B05213;
  assign memory[ 250] = 32'h06402CA3;
  assign memory[ 251] = 32'h07E05293;
  assign memory[ 252] = 32'h005024A3;
  assign memory[ 253] = 32'h20502AA3;
  assign memory[ 254] = 32'h0F605313;
  assign memory[ 255] = 32'h22602CA3;
  assign memory[ 256] = 32'h0F705393;
  assign memory[ 257] = 32'h24702423;
  assign memory[ 258] = 32'h0F805413;
  assign memory[ 259] = 32'h00802FA3;
  assign memory[ 260] = 32'h24802C23;
  assign memory[ 261] = 32'h0F905493;
  assign memory[ 262] = 32'h02902D23;
  assign memory[ 263] = 32'h2A9023A3;
  assign memory[ 264] = 32'h0FA05513;
  assign memory[ 265] = 32'h08A024A3;
  assign memory[ 266] = 32'h0FE05593;
  assign memory[ 267] = 32'h00B02523;
  assign memory[ 268] = 32'h20B02B23;
  assign memory[ 269] = 32'h1F405613;
  assign memory[ 270] = 32'h22C02723;
  assign memory[ 271] = 32'h1F505693;
  assign memory[ 272] = 32'h22D02D23;
  assign memory[ 273] = 32'h1F605713;
  assign memory[ 274] = 32'h02E02623;
  assign memory[ 275] = 32'h26E02423;
  assign memory[ 276] = 32'h1F705793;
  assign memory[ 277] = 32'h04F02523;
  assign memory[ 278] = 32'h2AF02BA3;
  assign memory[ 279] = 32'h1F805813;
  assign memory[ 280] = 32'h09002CA3;
  assign memory[ 281] = 32'h2D0023A3;
  assign memory[ 282] = 32'h1F905893;
  assign memory[ 283] = 32'h0B1024A3;
  assign memory[ 284] = 32'h2D102BA3;
  assign memory[ 285] = 32'h1FA05913;
  assign memory[ 286] = 32'h0B202CA3;
  assign memory[ 287] = 32'h2F2023A3;
  assign memory[ 288] = 32'h1FE05993;
  assign memory[ 289] = 32'h013025A3;
  assign memory[ 290] = 32'h21302BA3;
  assign memory[ 291] = 32'h3F605A13;
  assign memory[ 292] = 32'h03402023;
  assign memory[ 293] = 32'h234027A3;
  assign memory[ 294] = 32'h3F705A93;
  assign memory[ 295] = 32'h03502DA3;
  assign memory[ 296] = 32'h255024A3;
  assign memory[ 297] = 32'h3F805B13;
  assign memory[ 298] = 32'h05602D23;
  assign memory[ 299] = 32'h25602CA3;
  assign memory[ 300] = 32'h3F905B93;
  assign memory[ 301] = 32'h0D7024A3;
  assign memory[ 302] = 32'h27702C23;
  assign memory[ 303] = 32'h3FA05C13;
  assign memory[ 304] = 32'h0D802CA3;
  assign memory[ 305] = 32'h31802B23;
  assign memory[ 306] = 32'h3FE05C93;
  assign memory[ 307] = 32'h21902C23;
  assign memory[ 308] = 32'h3FF05D13;
  assign memory[ 309] = 32'h4BA02123;
  assign memory[ 310] = 32'h7F605D93;
  assign memory[ 311] = 32'h03B026A3;
  assign memory[ 312] = 32'h23B02DA3;
  assign memory[ 313] = 32'h7F705E13;
  assign memory[ 314] = 32'h07C02523;
  assign memory[ 315] = 32'h29C02423;
  assign memory[ 316] = 32'h7F805E93;
  assign memory[ 317] = 32'h0FD024A3;
  assign memory[ 318] = 32'h29D02C23;
  assign memory[ 319] = 32'h7F905093;
  assign memory[ 320] = 32'h10102423;
  assign memory[ 321] = 32'h2E102BA3;
  assign memory[ 322] = 32'h7FE05113;
  assign memory[ 323] = 32'h20202CA3;
  assign memory[ 324] = 32'h7FF05193;
  assign memory[ 325] = 32'h4A3020A3;
  assign memory[ 326] = 32'h7FB0D213;
  assign memory[ 327] = 32'h02402E23;
  assign memory[ 328] = 32'h22402823;
  assign memory[ 329] = 32'h7FC0D293;
  assign memory[ 330] = 32'h045025A3;
  assign memory[ 331] = 32'h22502E23;
  assign memory[ 332] = 32'h7FD0D313;
  assign memory[ 333] = 32'h06602D23;
  assign memory[ 334] = 32'h24602523;
  assign memory[ 335] = 32'h7FE0D393;
  assign memory[ 336] = 32'h08702523;
  assign memory[ 337] = 32'h24702D23;
  assign memory[ 338] = 32'h7FC15413;
  assign memory[ 339] = 32'h4A802023;
  assign memory[ 340] = 32'h00305F13;
  assign memory[ 341] = 32'h00B05F93;
  assign memory[ 342] = 32'h01FF1F33;
  assign memory[ 343] = 32'h7D505F93;
  assign memory[ 344] = 32'h01FF64B3;
  assign memory[ 345] = 32'h48902FA3;
  assign memory[ 346] = 32'h00605F13;
  assign memory[ 347] = 32'h00B05F93;
  assign memory[ 348] = 32'h01FF1F33;
  assign memory[ 349] = 32'h24405F93;
  assign memory[ 350] = 32'h01FF6533;
  assign memory[ 351] = 32'h4AA02823;
  assign memory[ 352] = 32'h5BC55F13;
  assign memory[ 353] = 32'h6B605F93;
  assign memory[ 354] = 32'h01FF65B3;
  assign memory[ 355] = 32'h48B02F23;
  assign memory[ 356] = 32'h12A5D613;
  assign memory[ 357] = 32'h30C023A3;
  assign memory[ 358] = 32'h00E05F13;
  assign memory[ 359] = 32'h00B05F93;
  assign memory[ 360] = 32'h01FF1F33;
  assign memory[ 361] = 32'h6B105F93;
  assign memory[ 362] = 32'h01FF66B3;
  assign memory[ 363] = 32'h48D02EA3;
  assign memory[ 364] = 32'h14F6DF13;
  assign memory[ 365] = 32'h7C005F93;
  assign memory[ 366] = 32'h01FF6733;
  assign memory[ 367] = 32'h08E02D23;
  assign memory[ 368] = 32'h00275793;
  assign memory[ 369] = 32'h24F025A3;
  assign memory[ 370] = 32'h00375813;
  assign memory[ 371] = 32'h31002BA3;
  assign memory[ 372] = 32'h01605F13;
  assign memory[ 373] = 32'h00B05F93;
  assign memory[ 374] = 32'h01FF1F33;
  assign memory[ 375] = 32'h50505F93;
  assign memory[ 376] = 32'h01FF68B3;
  assign memory[ 377] = 32'h4B102723;
  assign memory[ 378] = 32'h01905F13;
  assign memory[ 379] = 32'h00B05F93;
  assign memory[ 380] = 32'h01FF1F33;
  assign memory[ 381] = 32'h10F05F93;
  assign memory[ 382] = 32'h01FF6933;
  assign memory[ 383] = 32'h49202E23;
  assign memory[ 384] = 32'h01F05F13;
  assign memory[ 385] = 32'h00B05F93;
  assign memory[ 386] = 32'h01FF1F33;
  assign memory[ 387] = 32'h78205F93;
  assign memory[ 388] = 32'h01FF69B3;
  assign memory[ 389] = 32'h033020A3;
  assign memory[ 390] = 32'h0019DA13;
  assign memory[ 391] = 32'h03402123;
  assign memory[ 392] = 32'h0029DA93;
  assign memory[ 393] = 32'h03502723;
  assign memory[ 394] = 32'h0039DB13;
  assign memory[ 395] = 32'h036027A3;
  assign memory[ 396] = 32'h0049DB93;
  assign memory[ 397] = 32'h03702823;
  assign memory[ 398] = 32'h0059DC13;
  assign memory[ 399] = 32'h038028A3;
  assign memory[ 400] = 32'h0069DC93;
  assign memory[ 401] = 32'h03902923;
  assign memory[ 402] = 32'h23902EA3;
  assign memory[ 403] = 32'h0079DD13;
  assign memory[ 404] = 32'h03A02EA3;
  assign memory[ 405] = 32'h23A02F23;
  assign memory[ 406] = 32'h0089DD93;
  assign memory[ 407] = 32'h03B02F23;
  assign memory[ 408] = 32'h23B02FA3;
  assign memory[ 409] = 32'h0099DE13;
  assign memory[ 410] = 32'h03C02FA3;
  assign memory[ 411] = 32'h25C02023;
  assign memory[ 412] = 32'h00A9DE93;
  assign memory[ 413] = 32'h05D02023;
  assign memory[ 414] = 32'h25D02623;
  assign memory[ 415] = 32'h00B9D093;
  assign memory[ 416] = 32'h041020A3;
  assign memory[ 417] = 32'h241026A3;
  assign memory[ 418] = 32'h0010D113;
  assign memory[ 419] = 32'h04202123;
  assign memory[ 420] = 32'h24202723;
  assign memory[ 421] = 32'h0020D193;
  assign memory[ 422] = 32'h04302623;
  assign memory[ 423] = 32'h243027A3;
  assign memory[ 424] = 32'h0030D213;
  assign memory[ 425] = 32'h044026A3;
  assign memory[ 426] = 32'h24402823;
  assign memory[ 427] = 32'h0040D293;
  assign memory[ 428] = 32'h04502723;
  assign memory[ 429] = 32'h24502DA3;
  assign memory[ 430] = 32'h0050D313;
  assign memory[ 431] = 32'h046027A3;
  assign memory[ 432] = 32'h24602E23;
  assign memory[ 433] = 32'h0060D393;
  assign memory[ 434] = 32'h04702823;
  assign memory[ 435] = 32'h24702EA3;
  assign memory[ 436] = 32'h0070D413;
  assign memory[ 437] = 32'h048028A3;
  assign memory[ 438] = 32'h24802F23;
  assign memory[ 439] = 32'h0080D493;
  assign memory[ 440] = 32'h04902923;
  assign memory[ 441] = 32'h24902FA3;
  assign memory[ 442] = 32'h0090D513;
  assign memory[ 443] = 32'h04A02DA3;
  assign memory[ 444] = 32'h26A02023;
  assign memory[ 445] = 32'h00A0D593;
  assign memory[ 446] = 32'h04B02E23;
  assign memory[ 447] = 32'h26B024A3;
  assign memory[ 448] = 32'h00B0D613;
  assign memory[ 449] = 32'h04C02EA3;
  assign memory[ 450] = 32'h26C02523;
  assign memory[ 451] = 32'h00C0D693;
  assign memory[ 452] = 32'h04D02F23;
  assign memory[ 453] = 32'h26D025A3;
  assign memory[ 454] = 32'h00D0D713;
  assign memory[ 455] = 32'h04E02FA3;
  assign memory[ 456] = 32'h26E02623;
  assign memory[ 457] = 32'h00E0D793;
  assign memory[ 458] = 32'h06F02023;
  assign memory[ 459] = 32'h26F026A3;
  assign memory[ 460] = 32'h00F0D813;
  assign memory[ 461] = 32'h070020A3;
  assign memory[ 462] = 32'h27002723;
  assign memory[ 463] = 32'h0100D893;
  assign memory[ 464] = 32'h07102123;
  assign memory[ 465] = 32'h271027A3;
  assign memory[ 466] = 32'h0110D913;
  assign memory[ 467] = 32'h072025A3;
  assign memory[ 468] = 32'h27202823;
  assign memory[ 469] = 32'h0120D993;
  assign memory[ 470] = 32'h07302623;
  assign memory[ 471] = 32'h27302CA3;
  assign memory[ 472] = 32'h0130DA13;
  assign memory[ 473] = 32'h074026A3;
  assign memory[ 474] = 32'h27402D23;
  assign memory[ 475] = 32'h0140DA93;
  assign memory[ 476] = 32'h07502723;
  assign memory[ 477] = 32'h27502DA3;
  assign memory[ 478] = 32'h0150DB13;
  assign memory[ 479] = 32'h076027A3;
  assign memory[ 480] = 32'h27602E23;
  assign memory[ 481] = 32'h0160DB93;
  assign memory[ 482] = 32'h07702823;
  assign memory[ 483] = 32'h27702EA3;
  assign memory[ 484] = 32'h0170DC13;
  assign memory[ 485] = 32'h078028A3;
  assign memory[ 486] = 32'h27802F23;
  assign memory[ 487] = 32'h0180DC93;
  assign memory[ 488] = 32'h07902923;
  assign memory[ 489] = 32'h27902FA3;
  assign memory[ 490] = 32'h0190DD13;
  assign memory[ 491] = 32'h07A02DA3;
  assign memory[ 492] = 32'h29A02023;
  assign memory[ 493] = 32'h01A0DD93;
  assign memory[ 494] = 32'h07B02E23;
  assign memory[ 495] = 32'h29B024A3;
  assign memory[ 496] = 32'h01B0DE13;
  assign memory[ 497] = 32'h07C02EA3;
  assign memory[ 498] = 32'h29C02523;
  assign memory[ 499] = 32'h01C0DE93;
  assign memory[ 500] = 32'h07D02F23;
  assign memory[ 501] = 32'h29D025A3;
  assign memory[ 502] = 32'h01D0D093;
  assign memory[ 503] = 32'h06102FA3;
  assign memory[ 504] = 32'h28102623;
  assign memory[ 505] = 32'h0010D113;
  assign memory[ 506] = 32'h08202023;
  assign memory[ 507] = 32'h282026A3;
  assign memory[ 508] = 32'h0020D193;
  assign memory[ 509] = 32'h083020A3;
  assign memory[ 510] = 32'h28302723;
  assign memory[ 511] = 32'h0030D213;
  assign memory[ 512] = 32'h08402123;
  assign memory[ 513] = 32'h284027A3;
  assign memory[ 514] = 32'h0040D293;
  assign memory[ 515] = 32'h085025A3;
  assign memory[ 516] = 32'h28502823;
  assign memory[ 517] = 32'h0050D313;
  assign memory[ 518] = 32'h08602623;
  assign memory[ 519] = 32'h28602CA3;
  assign memory[ 520] = 32'h0060D393;
  assign memory[ 521] = 32'h087026A3;
  assign memory[ 522] = 32'h28702D23;
  assign memory[ 523] = 32'h0070D413;
  assign memory[ 524] = 32'h08802723;
  assign memory[ 525] = 32'h28802DA3;
  assign memory[ 526] = 32'h0080D493;
  assign memory[ 527] = 32'h089027A3;
  assign memory[ 528] = 32'h28902E23;
  assign memory[ 529] = 32'h0090D513;
  assign memory[ 530] = 32'h08A02823;
  assign memory[ 531] = 32'h28A02EA3;
  assign memory[ 532] = 32'h00A0D593;
  assign memory[ 533] = 32'h08B028A3;
  assign memory[ 534] = 32'h28B02F23;
  assign memory[ 535] = 32'h00B0D613;
  assign memory[ 536] = 32'h08C02923;
  assign memory[ 537] = 32'h28C02FA3;
  assign memory[ 538] = 32'h00C0D693;
  assign memory[ 539] = 32'h08D02DA3;
  assign memory[ 540] = 32'h2AD02023;
  assign memory[ 541] = 32'h00D0D713;
  assign memory[ 542] = 32'h08E02E23;
  assign memory[ 543] = 32'h2AE02423;
  assign memory[ 544] = 32'h00E0D793;
  assign memory[ 545] = 32'h08F02EA3;
  assign memory[ 546] = 32'h2AF024A3;
  assign memory[ 547] = 32'h00F0D813;
  assign memory[ 548] = 32'h09002F23;
  assign memory[ 549] = 32'h2B002523;
  assign memory[ 550] = 32'h0100D893;
  assign memory[ 551] = 32'h09102FA3;
  assign memory[ 552] = 32'h2B1025A3;
  assign memory[ 553] = 32'h0110D913;
  assign memory[ 554] = 32'h0B202023;
  assign memory[ 555] = 32'h2B202623;
  assign memory[ 556] = 32'h0120D993;
  assign memory[ 557] = 32'h0B3020A3;
  assign memory[ 558] = 32'h2B3026A3;
  assign memory[ 559] = 32'h0130DA13;
  assign memory[ 560] = 32'h0B402123;
  assign memory[ 561] = 32'h2B402723;
  assign memory[ 562] = 32'h0140DA93;
  assign memory[ 563] = 32'h0B502523;
  assign memory[ 564] = 32'h2B5027A3;
  assign memory[ 565] = 32'h0150DB13;
  assign memory[ 566] = 32'h0B6025A3;
  assign memory[ 567] = 32'h2B602823;
  assign memory[ 568] = 32'h0160DB93;
  assign memory[ 569] = 32'h0B702623;
  assign memory[ 570] = 32'h2B702C23;
  assign memory[ 571] = 32'h0170DC13;
  assign memory[ 572] = 32'h0B8026A3;
  assign memory[ 573] = 32'h2B802CA3;
  assign memory[ 574] = 32'h0180DC93;
  assign memory[ 575] = 32'h0B902723;
  assign memory[ 576] = 32'h2B902D23;
  assign memory[ 577] = 32'h0190DD13;
  assign memory[ 578] = 32'h0BA027A3;
  assign memory[ 579] = 32'h2BA02DA3;
  assign memory[ 580] = 32'h01A0DD93;
  assign memory[ 581] = 32'h0BB02823;
  assign memory[ 582] = 32'h2BB02E23;
  assign memory[ 583] = 32'h01B0DE13;
  assign memory[ 584] = 32'h0BC028A3;
  assign memory[ 585] = 32'h2BC02EA3;
  assign memory[ 586] = 32'h01C0DE93;
  assign memory[ 587] = 32'h0BD02923;
  assign memory[ 588] = 32'h2BD02F23;
  assign memory[ 589] = 32'h01D0D093;
  assign memory[ 590] = 32'h0A102D23;
  assign memory[ 591] = 32'h2A102FA3;
  assign memory[ 592] = 32'h0010D113;
  assign memory[ 593] = 32'h0A202DA3;
  assign memory[ 594] = 32'h2C202023;
  assign memory[ 595] = 32'h0020D193;
  assign memory[ 596] = 32'h0A302E23;
  assign memory[ 597] = 32'h2C302423;
  assign memory[ 598] = 32'h0030D213;
  assign memory[ 599] = 32'h0A402EA3;
  assign memory[ 600] = 32'h2C4024A3;
  assign memory[ 601] = 32'h0040D293;
  assign memory[ 602] = 32'h0A502F23;
  assign memory[ 603] = 32'h2C502523;
  assign memory[ 604] = 32'h0050D313;
  assign memory[ 605] = 32'h0A602FA3;
  assign memory[ 606] = 32'h2C6025A3;
  assign memory[ 607] = 32'h0060D393;
  assign memory[ 608] = 32'h0C702023;
  assign memory[ 609] = 32'h2C702623;
  assign memory[ 610] = 32'h0070D413;
  assign memory[ 611] = 32'h0C8020A3;
  assign memory[ 612] = 32'h2C8026A3;
  assign memory[ 613] = 32'h0080D493;
  assign memory[ 614] = 32'h0C902123;
  assign memory[ 615] = 32'h2C902723;
  assign memory[ 616] = 32'h0090D513;
  assign memory[ 617] = 32'h0CA02523;
  assign memory[ 618] = 32'h2CA027A3;
  assign memory[ 619] = 32'h00A0D593;
  assign memory[ 620] = 32'h0CB025A3;
  assign memory[ 621] = 32'h2CB02823;
  assign memory[ 622] = 32'h00B0D613;
  assign memory[ 623] = 32'h0CC02623;
  assign memory[ 624] = 32'h2CC02C23;
  assign memory[ 625] = 32'h00C0D693;
  assign memory[ 626] = 32'h0CD026A3;
  assign memory[ 627] = 32'h2CD02CA3;
  assign memory[ 628] = 32'h00D0D713;
  assign memory[ 629] = 32'h0CE02723;
  assign memory[ 630] = 32'h2CE02D23;
  assign memory[ 631] = 32'h00E0D793;
  assign memory[ 632] = 32'h0CF027A3;
  assign memory[ 633] = 32'h2CF02DA3;
  assign memory[ 634] = 32'h00F0D813;
  assign memory[ 635] = 32'h0D002823;
  assign memory[ 636] = 32'h2D002E23;
  assign memory[ 637] = 32'h0100D893;
  assign memory[ 638] = 32'h0D1028A3;
  assign memory[ 639] = 32'h2D102EA3;
  assign memory[ 640] = 32'h0110D913;
  assign memory[ 641] = 32'h0D202923;
  assign memory[ 642] = 32'h2D202F23;
  assign memory[ 643] = 32'h0120D993;
  assign memory[ 644] = 32'h0D302D23;
  assign memory[ 645] = 32'h2D302FA3;
  assign memory[ 646] = 32'h0130DA13;
  assign memory[ 647] = 32'h0D402DA3;
  assign memory[ 648] = 32'h2F402023;
  assign memory[ 649] = 32'h0140DA93;
  assign memory[ 650] = 32'h0D502E23;
  assign memory[ 651] = 32'h2F502423;
  assign memory[ 652] = 32'h0150DB13;
  assign memory[ 653] = 32'h0D602EA3;
  assign memory[ 654] = 32'h2F6024A3;
  assign memory[ 655] = 32'h0160DB93;
  assign memory[ 656] = 32'h0D702F23;
  assign memory[ 657] = 32'h2F702523;
  assign memory[ 658] = 32'h0170DC13;
  assign memory[ 659] = 32'h0D802FA3;
  assign memory[ 660] = 32'h2F8025A3;
  assign memory[ 661] = 32'h0180DC93;
  assign memory[ 662] = 32'h0F902023;
  assign memory[ 663] = 32'h2F902623;
  assign memory[ 664] = 32'h0190DD13;
  assign memory[ 665] = 32'h0FA020A3;
  assign memory[ 666] = 32'h2FA026A3;
  assign memory[ 667] = 32'h01A0DD93;
  assign memory[ 668] = 32'h0FB02123;
  assign memory[ 669] = 32'h2FB02723;
  assign memory[ 670] = 32'h01B0DE13;
  assign memory[ 671] = 32'h0FC02523;
  assign memory[ 672] = 32'h2FC027A3;
  assign memory[ 673] = 32'h01C0DE93;
  assign memory[ 674] = 32'h0FD025A3;
  assign memory[ 675] = 32'h2FD02823;
  assign memory[ 676] = 32'h01D0D093;
  assign memory[ 677] = 32'h0E102623;
  assign memory[ 678] = 32'h2E102C23;
  assign memory[ 679] = 32'h0010D113;
  assign memory[ 680] = 32'h0E2026A3;
  assign memory[ 681] = 32'h2E202CA3;
  assign memory[ 682] = 32'h0020D193;
  assign memory[ 683] = 32'h0E302723;
  assign memory[ 684] = 32'h2E302D23;
  assign memory[ 685] = 32'h0030D213;
  assign memory[ 686] = 32'h0E4027A3;
  assign memory[ 687] = 32'h2E402DA3;
  assign memory[ 688] = 32'h0040D293;
  assign memory[ 689] = 32'h0E502823;
  assign memory[ 690] = 32'h2E502E23;
  assign memory[ 691] = 32'h0050D313;
  assign memory[ 692] = 32'h0E6028A3;
  assign memory[ 693] = 32'h2E602EA3;
  assign memory[ 694] = 32'h0060D393;
  assign memory[ 695] = 32'h0E702923;
  assign memory[ 696] = 32'h2E702F23;
  assign memory[ 697] = 32'h0070D413;
  assign memory[ 698] = 32'h0E802CA3;
  assign memory[ 699] = 32'h2E802FA3;
  assign memory[ 700] = 32'h0080D493;
  assign memory[ 701] = 32'h0E902D23;
  assign memory[ 702] = 32'h30902023;
  assign memory[ 703] = 32'h0090D513;
  assign memory[ 704] = 32'h0EA02DA3;
  assign memory[ 705] = 32'h30A02423;
  assign memory[ 706] = 32'h00A0D593;
  assign memory[ 707] = 32'h0EB02E23;
  assign memory[ 708] = 32'h30B024A3;
  assign memory[ 709] = 32'h00B0D613;
  assign memory[ 710] = 32'h0EC02EA3;
  assign memory[ 711] = 32'h30C02523;
  assign memory[ 712] = 32'h00C0D693;
  assign memory[ 713] = 32'h0ED02F23;
  assign memory[ 714] = 32'h30D025A3;
  assign memory[ 715] = 32'h00D0D713;
  assign memory[ 716] = 32'h0EE02FA3;
  assign memory[ 717] = 32'h30E02623;
  assign memory[ 718] = 32'h00E0D793;
  assign memory[ 719] = 32'h10F02023;
  assign memory[ 720] = 32'h30F026A3;
  assign memory[ 721] = 32'h00F0D813;
  assign memory[ 722] = 32'h110020A3;
  assign memory[ 723] = 32'h31002723;
  assign memory[ 724] = 32'h0100D893;
  assign memory[ 725] = 32'h11102123;
  assign memory[ 726] = 32'h311027A3;
  assign memory[ 727] = 32'h0110D913;
  assign memory[ 728] = 32'h112024A3;
  assign memory[ 729] = 32'h31202823;
  assign memory[ 730] = 32'h0120D993;
  assign memory[ 731] = 32'h11302523;
  assign memory[ 732] = 32'h31302C23;
  assign memory[ 733] = 32'h0130DA13;
  assign memory[ 734] = 32'h114025A3;
  assign memory[ 735] = 32'h31402CA3;
  assign memory[ 736] = 32'h0140DA93;
  assign memory[ 737] = 32'h11502623;
  assign memory[ 738] = 32'h31502D23;
  assign memory[ 739] = 32'h0150DB13;
  assign memory[ 740] = 32'h116026A3;
  assign memory[ 741] = 32'h31602DA3;
  assign memory[ 742] = 32'h0160DB93;
  assign memory[ 743] = 32'h11702723;
  assign memory[ 744] = 32'h31702E23;
  assign memory[ 745] = 32'h0170DC13;
  assign memory[ 746] = 32'h118027A3;
  assign memory[ 747] = 32'h31802EA3;
  assign memory[ 748] = 32'h0180DC93;
  assign memory[ 749] = 32'h11902823;
  assign memory[ 750] = 32'h31902F23;
  assign memory[ 751] = 32'h0190DD13;
  assign memory[ 752] = 32'h11A028A3;
  assign memory[ 753] = 32'h31A02FA3;
  assign memory[ 754] = 32'h01A0DD93;
  assign memory[ 755] = 32'h11B02923;
  assign memory[ 756] = 32'h33B02023;
  assign memory[ 757] = 32'h01C0DE13;
  assign memory[ 758] = 32'h4BC027A3;
  assign memory[ 759] = 32'h01605F93;
  assign memory[ 760] = 32'h03205E93;
  assign memory[ 761] = 32'h01FE9EB3;
  assign memory[ 762] = 32'h00B05F93;
  assign memory[ 763] = 32'h16805F13;
  assign memory[ 764] = 32'h01FF1F33;
  assign memory[ 765] = 32'h01DF6EB3;
  assign memory[ 766] = 32'h39505F93;
  assign memory[ 767] = 32'h01DFEEB3;
  assign memory[ 768] = 32'h4BD02D23;
  assign memory[ 769] = 32'h01605F93;
  assign memory[ 770] = 32'h08305E93;
  assign memory[ 771] = 32'h01FE9EB3;
  assign memory[ 772] = 32'h00B05F93;
  assign memory[ 773] = 32'h4AC05F13;
  assign memory[ 774] = 32'h01FF1F33;
  assign memory[ 775] = 32'h01DF6EB3;
  assign memory[ 776] = 32'h04105F93;
  assign memory[ 777] = 32'h01DFE0B3;
  assign memory[ 778] = 32'h4A102C23;
  assign memory[ 779] = 32'h01605F93;
  assign memory[ 780] = 32'h0E005E93;
  assign memory[ 781] = 32'h01FE9EB3;
  assign memory[ 782] = 32'h00B05F93;
  assign memory[ 783] = 32'h62405F13;
  assign memory[ 784] = 32'h01FF1F33;
  assign memory[ 785] = 32'h01DF6EB3;
  assign memory[ 786] = 32'h6E905F93;
  assign memory[ 787] = 32'h01DFE133;
  assign memory[ 788] = 32'h4A202EA3;
  assign memory[ 789] = 32'h01605F93;
  assign memory[ 790] = 32'h12005E93;
  assign memory[ 791] = 32'h01FE9EB3;
  assign memory[ 792] = 32'h00B05F93;
  assign memory[ 793] = 32'h62405F13;
  assign memory[ 794] = 32'h01FF1F33;
  assign memory[ 795] = 32'h01DF6EB3;
  assign memory[ 796] = 32'h6E905F93;
  assign memory[ 797] = 32'h01DFE1B3;
  assign memory[ 798] = 32'h4A302CA3;
  assign memory[ 799] = 32'h06405F13;
  assign memory[ 800] = 32'h00B05F93;
  assign memory[ 801] = 32'h01FF1F33;
  assign memory[ 802] = 32'h7D005F93;
  assign memory[ 803] = 32'h01FF6A33;
  assign memory[ 804] = 32'h7D005A93;
  assign memory[ 805] = 32'h000A2E03;
  assign memory[ 806] = 32'h001A2E83;
  assign memory[ 807] = 32'h4BC021A3;
  assign memory[ 808] = 32'h4BD02223;
  assign memory[ 809] = 32'h00405093;
  assign memory[ 810] = 32'h401E5E33;
  assign memory[ 811] = 32'h401EDDB3;
  assign memory[ 812] = 32'h4BC022A3;
  assign memory[ 813] = 32'h4BB02323;
  assign memory[ 814] = 32'h00005093;
  assign memory[ 815] = 32'h00005113;
  assign memory[ 816] = 32'h00005193;
  assign memory[ 817] = 32'h00005213;
  assign memory[ 818] = 32'h00005293;
  assign memory[ 819] = 32'h00005313;
  assign memory[ 820] = 32'h01005D13;
  assign memory[ 821] = 32'h00805C93;
  assign memory[ 822] = 32'h00205C13;
  assign memory[ 823] = 32'h15C10063;
  assign memory[ 824] = 32'h03DD0533;
  assign memory[ 825] = 32'h02250533;
  assign memory[ 826] = 32'h00255513;
  assign memory[ 827] = 32'h13B08263;
  assign memory[ 828] = 32'h021D05B3;
  assign memory[ 829] = 32'h00A585B3;
  assign memory[ 830] = 32'h11820663;
  assign memory[ 831] = 32'h03DC8633;
  assign memory[ 832] = 32'h02460633;
  assign memory[ 833] = 32'h00B60633;
  assign memory[ 834] = 32'h0F818863;
  assign memory[ 835] = 32'h023C86B3;
  assign memory[ 836] = 32'h00C686B3;
  assign memory[ 837] = 32'h0D928C63;
  assign memory[ 838] = 32'h00D28733;
  assign memory[ 839] = 32'h0D930263;
  assign memory[ 840] = 32'h026E87B3;
  assign memory[ 841] = 32'h00E787B3;
  assign memory[ 842] = 32'h00FA07B3;
  assign memory[ 843] = 32'h0FF05993;
  assign memory[ 844] = 32'h0007A803;
  assign memory[ 845] = 32'h41A85833;
  assign memory[ 846] = 32'h01387833;
  assign memory[ 847] = 32'h0007A883;
  assign memory[ 848] = 32'h4198D8B3;
  assign memory[ 849] = 32'h0138F8B3;
  assign memory[ 850] = 32'h0007A903;
  assign memory[ 851] = 32'h01397933;
  assign memory[ 852] = 32'h4B802983;
  assign memory[ 853] = 32'h030999B3;
  assign memory[ 854] = 32'h4B902F03;
  assign memory[ 855] = 32'h031F1F33;
  assign memory[ 856] = 32'h01E989B3;
  assign memory[ 857] = 32'h4BA02F03;
  assign memory[ 858] = 32'h032F1F33;
  assign memory[ 859] = 32'h01E989B3;
  assign memory[ 860] = 32'h0109D993;
  assign memory[ 861] = 32'h0009DB13;
  assign memory[ 862] = 32'h4BB02983;
  assign memory[ 863] = 32'h030999B3;
  assign memory[ 864] = 32'h4BC02F03;
  assign memory[ 865] = 32'h031F1F33;
  assign memory[ 866] = 32'h01E989B3;
  assign memory[ 867] = 32'h4BD02F03;
  assign memory[ 868] = 32'h032F1F33;
  assign memory[ 869] = 32'h01E989B3;
  assign memory[ 870] = 32'h0809D993;
  assign memory[ 871] = 32'h019999B3;
  assign memory[ 872] = 32'h01698B33;
  assign memory[ 873] = 32'h4BE02983;
  assign memory[ 874] = 32'h031999B3;
  assign memory[ 875] = 32'h4BD02F03;
  assign memory[ 876] = 32'h030F1F33;
  assign memory[ 877] = 32'h01E989B3;
  assign memory[ 878] = 32'h4BF02F03;
  assign memory[ 879] = 32'h032F1F33;
  assign memory[ 880] = 32'h01E989B3;
  assign memory[ 881] = 32'h0809D993;
  assign memory[ 882] = 32'h01A999B3;
  assign memory[ 883] = 32'h01698B33;
  assign memory[ 884] = 32'h016AA023;
  assign memory[ 885] = 32'h001ADA93;
  assign memory[ 886] = 32'h00135313;
  assign memory[ 887] = 32'hF40000E3;
  assign memory[ 888] = 32'h00005313;
  assign memory[ 889] = 32'h0012D293;
  assign memory[ 890] = 32'hF20006E3;
  assign memory[ 891] = 32'h00005293;
  assign memory[ 892] = 32'h0011D193;
  assign memory[ 893] = 32'hF0000AE3;
  assign memory[ 894] = 32'h00005193;
  assign memory[ 895] = 32'h00125213;
  assign memory[ 896] = 32'hEE000CE3;
  assign memory[ 897] = 32'h00005213;
  assign memory[ 898] = 32'h0010D093;
  assign memory[ 899] = 32'hEE0000E3;
  assign memory[ 900] = 32'h00005093;
  assign memory[ 901] = 32'h00115113;
  assign memory[ 902] = 32'hEC0002E3;
  assign memory[ 903] = 32'h06405F13;
  assign memory[ 904] = 32'h00B05F93;
  assign memory[ 905] = 32'h01FF1F33;
  assign memory[ 906] = 32'h7D005F93;
  assign memory[ 907] = 32'h01FF6533;
  assign memory[ 908] = 32'h06505F13;
  assign memory[ 909] = 32'h00B05F93;
  assign memory[ 910] = 32'h01FF1F33;
  assign memory[ 911] = 32'h3D205F93;
  assign memory[ 912] = 32'h01FF65B3;
  assign memory[ 913] = 32'h00B50863;
  assign memory[ 914] = 32'h00052023;
  assign memory[ 915] = 32'h00155513;
  assign memory[ 916] = 32'hFE000AE3;
  assign memory[ 917] = 32'h02005D13;
  assign memory[ 918] = 32'h06405F13;
  assign memory[ 919] = 32'h00B05F93;
  assign memory[ 920] = 32'h01FF1F33;
  assign memory[ 921] = 32'h7D005F93;
  assign memory[ 922] = 32'h01FF6CB3;
  assign memory[ 923] = 32'h5E000663;
  assign memory[ 924] = 32'h00005093;
  assign memory[ 925] = 32'h04005113;
  assign memory[ 926] = 32'h00208E63;
  assign memory[ 927] = 32'h5800A183;
  assign memory[ 928] = 32'hF801D193;
  assign memory[ 929] = 32'h5C30A023;
  assign memory[ 930] = 32'h5800A023;
  assign memory[ 931] = 32'h0010D093;
  assign memory[ 932] = 32'hFE0004E3;
  assign memory[ 933] = 32'h14000C63;
  assign memory[ 934] = 32'h00005413;
  assign memory[ 935] = 32'h06405F13;
  assign memory[ 936] = 32'h00B05F93;
  assign memory[ 937] = 32'h01FF1F33;
  assign memory[ 938] = 32'h43F05F93;
  assign memory[ 939] = 32'h01FF6A33;
  assign memory[ 940] = 32'hF3605F13;
  assign memory[ 941] = 32'h00B05F93;
  assign memory[ 942] = 32'h01FF1F33;
  assign memory[ 943] = 32'h78105F93;
  assign memory[ 944] = 32'h01FF6AB3;
  assign memory[ 945] = 32'h03205F13;
  assign memory[ 946] = 32'h00B05F93;
  assign memory[ 947] = 32'h01FF1F33;
  assign memory[ 948] = 32'h22005F93;
  assign memory[ 949] = 32'h01FF6B33;
  assign memory[ 950] = 32'h009A5663;
  assign memory[ 951] = 32'h015484B3;
  assign memory[ 952] = 32'hFE000CE3;
  assign memory[ 953] = 32'h009B5C63;
  assign memory[ 954] = 32'h00105413;
  assign memory[ 955] = 32'hFFFA6A13;
  assign memory[ 956] = 32'h001A5A13;
  assign memory[ 957] = 32'h014484B3;
  assign memory[ 958] = 32'h00000C63;
  assign memory[ 959] = 32'hFFFB6B13;
  assign memory[ 960] = 32'h001B5B13;
  assign memory[ 961] = 32'h0164D663;
  assign memory[ 962] = 32'h00105413;
  assign memory[ 963] = 32'h014484B3;
  assign memory[ 964] = 32'h00005513;
  assign memory[ 965] = 32'h4A0023A3;
  assign memory[ 966] = 32'h4A002423;
  assign memory[ 967] = 32'h4A0024A3;
  assign memory[ 968] = 32'h4A002523;
  assign memory[ 969] = 32'h4A0025A3;
  assign memory[ 970] = 32'h4A002623;
  assign memory[ 971] = 32'h4A0026A3;
  assign memory[ 972] = 32'h00005393;
  assign memory[ 973] = 32'h00705B13;
  assign memory[ 974] = 32'h03638C63;
  assign memory[ 975] = 32'h02A4D063;
  assign memory[ 976] = 32'h49C3AA03;
  assign memory[ 977] = 32'hFFFA6A13;
  assign memory[ 978] = 32'h001A5A13;
  assign memory[ 979] = 32'h01450533;
  assign memory[ 980] = 32'h00105A93;
  assign memory[ 981] = 32'h4B53A3A3;
  assign memory[ 982] = 32'h00000863;
  assign memory[ 983] = 32'h49C3AA03;
  assign memory[ 984] = 32'h01450533;
  assign memory[ 985] = 32'h4A03A3A3;
  assign memory[ 986] = 32'h0013D393;
  assign memory[ 987] = 32'hFC0006E3;
  assign memory[ 988] = 32'h01305F13;
  assign memory[ 989] = 32'h00B05F93;
  assign memory[ 990] = 32'h01FF1F33;
  assign memory[ 991] = 32'h37505F93;
  assign memory[ 992] = 32'h01FF60B3;
  assign memory[ 993] = 32'h00005113;
  assign memory[ 994] = 32'h00605393;
  assign memory[ 995] = 32'h00105A93;
  assign memory[ 996] = 32'hFFF05B93;
  assign memory[ 997] = 32'h05738063;
  assign memory[ 998] = 32'h4A73AA03;
  assign memory[ 999] = 32'h40715B33;
  assign memory[1000] = 32'h015A1C63;
  assign memory[1001] = 32'hFFFB6B13;
  assign memory[1002] = 32'h001B5B13;
  assign memory[1003] = 32'h016080B3;
  assign memory[1004] = 32'h4070DB33;
  assign memory[1005] = 32'h00000A63;
  assign memory[1006] = 32'h016080B3;
  assign memory[1007] = 32'h4070DB33;
  assign memory[1008] = 32'hFFFB6B13;
  assign memory[1009] = 32'h001B5B13;
  assign memory[1010] = 32'h002B0133;
  assign memory[1011] = 32'hFFF3D393;
  assign memory[1012] = 32'hFC0002E3;
  assign memory[1013] = 32'h01541663;
  assign memory[1014] = 32'hFFF0E093;
  assign memory[1015] = 32'h0010D093;
  assign memory[1016] = 32'h00105A93;
  assign memory[1017] = 32'h060C0E63;
  assign memory[1018] = 32'h095C0E63;
  assign memory[1019] = 32'h00805793;
  assign memory[1020] = 32'h00205893;
  assign memory[1021] = 32'h00005193;
  assign memory[1022] = 32'h00005213;
  assign memory[1023] = 32'h00005293;
  assign memory[1024] = 32'h00005313;
  assign memory[1025] = 32'h10F18E63;
  assign memory[1026] = 32'h00019663;
  assign memory[1027] = 32'h4AE02583;
  assign memory[1028] = 32'h00000463;
  assign memory[1029] = 32'h4AF02583;
  assign memory[1030] = 32'h0EF20E63;
  assign memory[1031] = 32'h00021663;
  assign memory[1032] = 32'h4AE02603;
  assign memory[1033] = 32'h00000463;
  assign memory[1034] = 32'h4AF02603;
  assign memory[1035] = 32'h00005713;
  assign memory[1036] = 32'h06F28A63;
  assign memory[1037] = 32'h06F30263;
  assign memory[1038] = 32'h02F28833;
  assign memory[1039] = 32'h00680833;
  assign memory[1040] = 32'h5C082683;
  assign memory[1041] = 32'h025884B3;
  assign memory[1042] = 32'h0014D493;
  assign memory[1043] = 32'h023484B3;
  assign memory[1044] = 32'h4B002B83;
  assign memory[1045] = 32'h037484B3;
  assign memory[1046] = 32'h00005C13;
  assign memory[1047] = 32'hE2000EE3;
  assign memory[1048] = 32'h021686B3;
  assign memory[1049] = 32'h40F6D6B3;
  assign memory[1050] = 32'h026884B3;
  assign memory[1051] = 32'h0014D493;
  assign memory[1052] = 32'h024484B3;
  assign memory[1053] = 32'h4B002B83;
  assign memory[1054] = 32'h037484B3;
  assign memory[1055] = 32'h00105C13;
  assign memory[1056] = 32'hE0000CE3;
  assign memory[1057] = 32'h021686B3;
  assign memory[1058] = 32'h40F6D6B3;
  assign memory[1059] = 32'h00D70733;
  assign memory[1060] = 32'h00135313;
  assign memory[1061] = 32'hFA0000E3;
  assign memory[1062] = 32'h00005313;
  assign memory[1063] = 32'h0012D293;
  assign memory[1064] = 32'hF80008E3;
  assign memory[1065] = 32'h02C59833;
  assign memory[1066] = 32'h02C586B3;
  assign memory[1067] = 32'h01605F93;
  assign memory[1068] = 32'h1FF05E93;
  assign memory[1069] = 32'h01FE9EB3;
  assign memory[1070] = 32'h00B05F93;
  assign memory[1071] = 32'h7FF05F13;
  assign memory[1072] = 32'h01FF1F33;
  assign memory[1073] = 32'h01DF6EB3;
  assign memory[1074] = 32'h7FF05F93;
  assign memory[1075] = 32'h01DFEAB3;
  assign memory[1076] = 32'h0156F6B3;
  assign memory[1077] = 32'h00F05913;
  assign memory[1078] = 32'h01281833;
  assign memory[1079] = 32'h00195913;
  assign memory[1080] = 32'h4126D6B3;
  assign memory[1081] = 32'h0106E6B3;
  assign memory[1082] = 32'h02E696B3;
  assign memory[1083] = 32'h00305913;
  assign memory[1084] = 32'h4126D6B3;
  assign memory[1085] = 32'h00068463;
  assign memory[1086] = 32'h0016D693;
  assign memory[1087] = 32'h02F18833;
  assign memory[1088] = 32'h01020833;
  assign memory[1089] = 32'h58D82023;
  assign memory[1090] = 32'h00005293;
  assign memory[1091] = 32'h00125213;
  assign memory[1092] = 32'hF00004E3;
  assign memory[1093] = 32'h00005213;
  assign memory[1094] = 32'h0011D193;
  assign memory[1095] = 32'hEE0004E3;
  assign memory[1096] = 32'h41C05113;
  assign memory[1097] = 32'h000E1463;
  assign memory[1098] = 32'h45C05113;
  assign memory[1099] = 32'h00005093;
  assign memory[1100] = 32'h04005293;
  assign memory[1101] = 32'h01005393;
  assign memory[1102] = 32'h02508463;
  assign memory[1103] = 32'h00208333;
  assign memory[1104] = 32'h00032183;
  assign memory[1105] = 32'h5800A203;
  assign memory[1106] = 32'h024181B3;
  assign memory[1107] = 32'h4071D1B3;
  assign memory[1108] = 32'h5800A023;
  assign memory[1109] = 32'h5C30A023;
  assign memory[1110] = 32'h0010D093;
  assign memory[1111] = 32'hFC000EE3;
  assign memory[1112] = 32'h00005093;
  assign memory[1113] = 32'h00005113;
  assign memory[1114] = 32'h00005293;
  assign memory[1115] = 32'h00105193;
  assign memory[1116] = 32'h00005213;
  assign memory[1117] = 32'h00705313;
  assign memory[1118] = 32'h00805393;
  assign memory[1119] = 32'h00105493;
  assign memory[1120] = 32'h4B4E2E83;
  assign memory[1121] = 32'h5C002D83;
  assign memory[1122] = 32'hFFFEEE93;
  assign memory[1123] = 32'h001EDE93;
  assign memory[1124] = 32'h01DD85B3;
  assign memory[1125] = 32'h4BBE2A23;
  assign memory[1126] = 32'h58B02023;
  assign memory[1127] = 32'h08001463;
  assign memory[1128] = 32'h00008663;
  assign memory[1129] = 32'h00608463;
  assign memory[1130] = 32'h00000863;
  assign memory[1131] = 32'h00115113;
  assign memory[1132] = 32'h00105213;
  assign memory[1133] = 32'h00000C63;
  assign memory[1134] = 32'h00010663;
  assign memory[1135] = 32'h00610463;
  assign memory[1136] = 32'h00000663;
  assign memory[1137] = 32'h0010D093;
  assign memory[1138] = 32'h00105213;
  assign memory[1139] = 32'h02921263;
  assign memory[1140] = 32'h00005213;
  assign memory[1141] = 32'hFFF1E193;
  assign memory[1142] = 32'h0011D193;
  assign memory[1143] = 32'h0012D293;
  assign memory[1144] = 32'h02710633;
  assign memory[1145] = 32'h00160633;
  assign memory[1146] = 32'h5C062583;
  assign memory[1147] = 32'h58B2A023;
  assign memory[1148] = 32'h00611663;
  assign memory[1149] = 32'h00609463;
  assign memory[1150] = 32'h02000663;
  assign memory[1151] = 32'h0012D293;
  assign memory[1152] = 32'hFFF1E693;
  assign memory[1153] = 32'h0016D693;
  assign memory[1154] = 32'h001680B3;
  assign memory[1155] = 32'h00310133;
  assign memory[1156] = 32'h02710633;
  assign memory[1157] = 32'h00160633;
  assign memory[1158] = 32'h5C062583;
  assign memory[1159] = 32'h58B2A023;
  assign memory[1160] = 32'hF6000EE3;
  assign memory[1161] = 32'h000E1C63;
  assign memory[1162] = 32'h00005513;
  assign memory[1163] = 32'h00C05593;
  assign memory[1164] = 32'h01805613;
  assign memory[1165] = 32'h11305693;
  assign memory[1166] = 32'h00000A63;
  assign memory[1167] = 32'h20E05513;
  assign memory[1168] = 32'h21A05593;
  assign memory[1169] = 32'h22605613;
  assign memory[1170] = 32'h32105693;
  assign memory[1171] = 32'h06000663;
  assign memory[1172] = 32'h00005713;
  assign memory[1173] = 32'h00005793;
  assign memory[1174] = 32'h00105893;
  assign memory[1175] = 32'h0000D863;
  assign memory[1176] = 32'hFFF0E093;
  assign memory[1177] = 32'h0010D093;
  assign memory[1178] = 32'h00105793;
  assign memory[1179] = 32'h0000D113;
  assign memory[1180] = 32'h00008863;
  assign memory[1181] = 32'h4110D0B3;
  assign memory[1182] = 32'h00175713;
  assign memory[1183] = 32'hFE000AE3;
  assign memory[1184] = 32'h00075193;
  assign memory[1185] = 32'h03179263;
  assign memory[1186] = 32'h00005813;
  assign memory[1187] = 32'h00070A63;
  assign memory[1188] = 32'h01181833;
  assign memory[1189] = 32'h00185813;
  assign memory[1190] = 32'hFFF75713;
  assign memory[1191] = 32'hFE0008E3;
  assign memory[1192] = 32'hFFF16113;
  assign memory[1193] = 32'h01017133;
  assign memory[1194] = 32'h00105993;
  assign memory[1195] = 32'h0A0C0E63;
  assign memory[1196] = 32'h133C0463;
  assign memory[1197] = 32'h9C0004E3;
  assign memory[1198] = 32'h0A000263;
  assign memory[1199] = 32'h000CA703;
  assign memory[1200] = 32'h025D4263;
  assign memory[1201] = 32'hFFF2E293;
  assign memory[1202] = 32'h0012D293;
  assign memory[1203] = 32'h005D0933;
  assign memory[1204] = 32'h01221933;
  assign memory[1205] = 32'h01270733;
  assign memory[1206] = 32'h00ECA023;
  assign memory[1207] = 32'h005D0D33;
  assign memory[1208] = 32'h04000E63;
  assign memory[1209] = 32'hFFFD6993;
  assign memory[1210] = 32'h0019D993;
  assign memory[1211] = 32'h01328933;
  assign memory[1212] = 32'h41225933;
  assign memory[1213] = 32'h01276733;
  assign memory[1214] = 32'h00ECA023;
  assign memory[1215] = 32'h013282B3;
  assign memory[1216] = 32'h0002D793;
  assign memory[1217] = 32'h00005813;
  assign memory[1218] = 32'h00105993;
  assign memory[1219] = 32'h00078A63;
  assign memory[1220] = 32'h01381833;
  assign memory[1221] = 32'h00185813;
  assign memory[1222] = 32'hFFF7D793;
  assign memory[1223] = 32'hFE0008E3;
  assign memory[1224] = 32'h00487833;
  assign memory[1225] = 32'hFFF2E993;
  assign memory[1226] = 32'h0019D993;
  assign memory[1227] = 32'h0209DD13;
  assign memory[1228] = 32'h01A818B3;
  assign memory[1229] = 32'h001CDC93;
  assign memory[1230] = 32'h011CA023;
  assign memory[1231] = 32'h00105993;
  assign memory[1232] = 32'h00205913;
  assign memory[1233] = 32'h00305293;
  assign memory[1234] = 32'h040B8263;
  assign memory[1235] = 32'h073B8E63;
  assign memory[1236] = 32'h0B2B8C63;
  assign memory[1237] = 32'h0C5B8A63;
  assign memory[1238] = 32'h920002E3;
  assign memory[1239] = 32'h58002083;
  assign memory[1240] = 32'h00005C13;
  assign memory[1241] = 32'hEE0006E3;
  assign memory[1242] = 32'h00350733;
  assign memory[1243] = 32'h00072303;
  assign memory[1244] = 32'h00358733;
  assign memory[1245] = 32'h00072383;
  assign memory[1246] = 32'h00331233;
  assign memory[1247] = 32'h00220233;
  assign memory[1248] = 32'h007182B3;
  assign memory[1249] = 32'h00005B93;
  assign memory[1250] = 32'hF2000AE3;
  assign memory[1251] = 32'h00005493;
  assign memory[1252] = 32'h00105A13;
  assign memory[1253] = 32'h04005A93;
  assign memory[1254] = 32'h00F05B13;
  assign memory[1255] = 32'h075A0C63;
  assign memory[1256] = 32'h580A2783;
  assign memory[1257] = 32'h00079663;
  assign memory[1258] = 32'h0014D493;
  assign memory[1259] = 32'h06000063;
  assign memory[1260] = 32'h009B5E63;
  assign memory[1261] = 32'hFF04D493;
  assign memory[1262] = 32'h0F062203;
  assign memory[1263] = 32'h0F06A283;
  assign memory[1264] = 32'h00105B93;
  assign memory[1265] = 32'hEE000CE3;
  assign memory[1266] = 32'hFE0004E3;
  assign memory[1267] = 32'h580A2083;
  assign memory[1268] = 32'h00105C13;
  assign memory[1269] = 32'hE6000EE3;
  assign memory[1270] = 32'h00405893;
  assign memory[1271] = 32'h01149433;
  assign memory[1272] = 32'h00340433;
  assign memory[1273] = 32'h00860733;
  assign memory[1274] = 32'h00072303;
  assign memory[1275] = 32'h00868733;
  assign memory[1276] = 32'h00072383;
  assign memory[1277] = 32'h00331233;
  assign memory[1278] = 32'h00220233;
  assign memory[1279] = 32'h007182B3;
  assign memory[1280] = 32'h00205B93;
  assign memory[1281] = 32'hEA000CE3;
  assign memory[1282] = 32'h00005493;
  assign memory[1283] = 32'h001A5A13;
  assign memory[1284] = 32'hF80006E3;
  assign memory[1285] = 32'h00048A63;
  assign memory[1286] = 32'h00062203;
  assign memory[1287] = 32'h0006A283;
  assign memory[1288] = 32'h00305B93;
  assign memory[1289] = 32'hE8000CE3;
  assign memory[1290] = 32'h0C805F13;
  assign memory[1291] = 32'h00B05F93;
  assign memory[1292] = 32'h01FF1F33;
  assign memory[1293] = 32'h7D005F93;
  assign memory[1294] = 32'h01FF6133;
  assign memory[1295] = 32'h01A12023;
  assign memory[1296] = 32'h00005093;
  assign memory[1297] = 32'h00105113;
  assign memory[1298] = 32'h00205193;
  assign memory[1299] = 32'h0C1E0463;
  assign memory[1300] = 32'h0E2E0E63;
  assign memory[1301] = 32'h123E0263;
  assign memory[1302] = 32'h4A0028A3;
  assign memory[1303] = 32'h4A002923;
  assign memory[1304] = 32'h4A0029A3;
  assign memory[1305] = 32'h4A002A23;
  assign memory[1306] = 32'h4A002AA3;
  assign memory[1307] = 32'h4A002B23;
  assign memory[1308] = 32'h10005093;
  assign memory[1309] = 32'h4A502103;
  assign memory[1310] = 32'h022080B3;
  assign memory[1311] = 32'h4A602103;
  assign memory[1312] = 32'h02208233;
  assign memory[1313] = 32'h4A402BA3;
  assign memory[1314] = 32'h00005093;
  assign memory[1315] = 32'h00005113;
  assign memory[1316] = 32'h00005193;
  assign memory[1317] = 32'h12408463;
  assign memory[1318] = 32'h7D00A303;
  assign memory[1319] = 32'h0FF05513;
  assign memory[1320] = 32'h00805593;
  assign memory[1321] = 32'h01005613;
  assign memory[1322] = 32'h00657333;
  assign memory[1323] = 32'h4C612023;
  assign memory[1324] = 32'h7D00A303;
  assign memory[1325] = 32'h40B35333;
  assign memory[1326] = 32'h00A37333;
  assign memory[1327] = 32'h50012383;
  assign memory[1328] = 32'h00730333;
  assign memory[1329] = 32'h50612023;
  assign memory[1330] = 32'h7D00A303;
  assign memory[1331] = 32'h54012383;
  assign memory[1332] = 32'h40C35333;
  assign memory[1333] = 32'h00A37333;
  assign memory[1334] = 32'h00730333;
  assign memory[1335] = 32'h54612023;
  assign memory[1336] = 32'h03F05313;
  assign memory[1337] = 32'h0C611663;
  assign memory[1338] = 32'h4A1028A3;
  assign memory[1339] = 32'h4A3029A3;
  assign memory[1340] = 32'h04005313;
  assign memory[1341] = 32'h00005393;
  assign memory[1342] = 32'h00638A63;
  assign memory[1343] = 32'h4C03A483;
  assign memory[1344] = 32'h5893A023;
  assign memory[1345] = 32'h0013D393;
  assign memory[1346] = 32'hFE0008E3;
  assign memory[1347] = 32'h00005E13;
  assign memory[1348] = 32'h960000E3;
  assign memory[1349] = 32'h4B302183;
  assign memory[1350] = 32'h00305413;
  assign memory[1351] = 32'h08819063;
  assign memory[1352] = 32'h04005313;
  assign memory[1353] = 32'h00005393;
  assign memory[1354] = 32'h00638E63;
  assign memory[1355] = 32'h5003A483;
  assign memory[1356] = 32'h00205293;
  assign memory[1357] = 32'h4054D4B3;
  assign memory[1358] = 32'h5893A023;
  assign memory[1359] = 32'h0013D393;
  assign memory[1360] = 32'hFE0004E3;
  assign memory[1361] = 32'h00105E13;
  assign memory[1362] = 32'h920004E3;
  assign memory[1363] = 32'h04005313;
  assign memory[1364] = 32'h00005393;
  assign memory[1365] = 32'h00638E63;
  assign memory[1366] = 32'h5403A483;
  assign memory[1367] = 32'h00205293;
  assign memory[1368] = 32'h4054D4B3;
  assign memory[1369] = 32'h5893A023;
  assign memory[1370] = 32'h0013D393;
  assign memory[1371] = 32'hFE0004E3;
  assign memory[1372] = 32'h00205E13;
  assign memory[1373] = 32'h8E000EE3;
  assign memory[1374] = 32'h04005313;
  assign memory[1375] = 32'h00005393;
  assign memory[1376] = 32'h00638A63;
  assign memory[1377] = 32'h5003A023;
  assign memory[1378] = 32'h5403A023;
  assign memory[1379] = 32'h0013D393;
  assign memory[1380] = 32'hFE0008E3;
  assign memory[1381] = 32'h00005193;
  assign memory[1382] = 32'h00000463;
  assign memory[1383] = 32'h0011D193;
  assign memory[1384] = 32'h00005113;
  assign memory[1385] = 32'h4B102083;
  assign memory[1386] = 32'h4B702203;
  assign memory[1387] = 32'h00000463;
  assign memory[1388] = 32'h00115113;
  assign memory[1389] = 32'h0010D093;
  assign memory[1390] = 32'hEC000EE3;
  assign memory[1391] = 32'h00005693;
  assign memory[1392] = 32'h00105093;
  assign memory[1393] = 32'h000D0A63;
  assign memory[1394] = 32'h001696B3;
  assign memory[1395] = 32'h0016D693;
  assign memory[1396] = 32'hFFFD5D13;
  assign memory[1397] = 32'hFE0008E3;
  assign memory[1398] = 32'h000CA103;
  assign memory[1399] = 32'h002686B3;
  assign memory[1400] = 32'h00DCA023;
  assign memory[1401] = 32'h00405F13;
  assign memory[1402] = 32'h00B05F93;
  assign memory[1403] = 32'h01FF1F33;
  assign memory[1404] = 32'h70F05F93;
  assign memory[1405] = 32'h01FF6FB3;

endmodule
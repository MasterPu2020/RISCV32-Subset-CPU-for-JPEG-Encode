//----------------------------------------------------------------
// JPEG encoding system on chip top module testbench
// Last Modified Date: 2023/7/17
// Version: 1.0
// Author: Clark Pu
//----------------------------------------------------------------

